library verilog;
use verilog.vl_types.all;
entity newfive_add_three_vlg_vec_tst is
end newfive_add_three_vlg_vec_tst;
