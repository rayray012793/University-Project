library verilog;
use verilog.vl_types.all;
entity newfulladder_vlg_vec_tst is
end newfulladder_vlg_vec_tst;
