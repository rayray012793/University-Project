library verilog;
use verilog.vl_types.all;
entity binarydowncounter_vlg_vec_tst is
end binarydowncounter_vlg_vec_tst;
