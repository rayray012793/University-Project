library verilog;
use verilog.vl_types.all;
entity binary_to_bcd_full_vlg_vec_tst is
end binary_to_bcd_full_vlg_vec_tst;
