library verilog;
use verilog.vl_types.all;
entity segementdecoder7_vlg_vec_tst is
end segementdecoder7_vlg_vec_tst;
