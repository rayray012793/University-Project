library verilog;
use verilog.vl_types.all;
entity binarytobcd_tb is
end binarytobcd_tb;
