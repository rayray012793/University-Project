library verilog;
use verilog.vl_types.all;
entity five_add_three_vlg_vec_tst is
end five_add_three_vlg_vec_tst;
