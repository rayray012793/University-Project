library verilog;
use verilog.vl_types.all;
entity binarytobcd_vlg_vec_tst is
end binarytobcd_vlg_vec_tst;
