library verilog;
use verilog.vl_types.all;
entity binaryupcounter_vlg_vec_tst is
end binaryupcounter_vlg_vec_tst;
