library verilog;
use verilog.vl_types.all;
entity segement7decoderverilog_vlg_check_tst is
    port(
        seg_out         : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end segement7decoderverilog_vlg_check_tst;
