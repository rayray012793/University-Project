library verilog;
use verilog.vl_types.all;
entity segement7decoderverilog_vlg_vec_tst is
end segement7decoderverilog_vlg_vec_tst;
