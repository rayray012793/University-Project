library verilog;
use verilog.vl_types.all;
entity new_binaryBCD_vlg_vec_tst is
end new_binaryBCD_vlg_vec_tst;
