library verilog;
use verilog.vl_types.all;
entity binaryupcounter_vlg_check_tst is
    port(
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        y3              : in     vl_logic;
        y4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end binaryupcounter_vlg_check_tst;
