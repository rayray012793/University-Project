library verilog;
use verilog.vl_types.all;
entity newfulladder_vlg_check_tst is
    port(
        C4              : in     vl_logic;
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        O3              : in     vl_logic;
        O4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end newfulladder_vlg_check_tst;
