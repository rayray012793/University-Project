library verilog;
use verilog.vl_types.all;
entity segementdecoder7 is
    port(
        a               : out    vl_logic;
        inputB          : in     vl_logic;
        inputD          : in     vl_logic;
        inputC          : in     vl_logic;
        inputA          : in     vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic
    );
end segementdecoder7;
